library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.all;

ENTITY DECODER IS --74_LS_42 MODIFICADO 
PORT (
	ENABLE_DEC: IN STD_LOGIC;
	IND: IN STD_LOGIC_VECTOR(7 downto 0);
	ADD,ADDC,CMP,INC,NOTT,MOVE,BZ,RETI: OUT STD_LOGIC;
	ST,LD,CLR,SHRR,SHLL,SUB,DEC,JMP: OUT STD_LOGIC;
	MODE: OUT STD_LOGIC;
	ADRS: OUT STD_LOGIC;
	OP1: OUT STD_LOGIC_VECTOR(2 downto 0);
	OP2: OUT STD_LOGIC_VECTOR (2 downto 0)
);
END DECODER;

ARCHITECTURE ESTRUCTURAL OF DECODER IS
BEGIN
PROCESS (ENABLE_DEC, IND)
    VARIABLE LECTURA: STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE MODO: STD_LOGIC;
BEGIN
    LECTURA := IND (7 DOWNTO 3);
    MODO := IND (2);
	IF LECTURA = "00000" THEN
	ADD <= '1';
	END IF;
	IF LECTURA = "00001" THEN
		ADDC <= '1';
	END IF;
	IF LECTURA = "00010" THEN
		CMP <= '1';
	END IF;
	IF LECTURA = "00011" THEN
		INC <= '1';
	END IF;
	IF LECTURA = "00100" THEN
		NOTT <= '1';
	END IF;
	IF LECTURA = "00110" THEN
		MOVE <= '1';
	END IF;
	IF LECTURA = "00111" THEN
		BZ <= '1';
	END IF;
	IF LECTURA = "01000" THEN
		RETI <= '1';
	END IF;
	IF LECTURA = "01011" THEN
		ST <= '1';
	END IF;
	IF LECTURA = "01100" THEN
		LD <= '1';
	END IF;
	IF LECTURA = "01101" THEN
		CLR <= '1';
	END IF;
	IF LECTURA = "01110" THEN
		SHRR <= '1';
	END IF;
	IF LECTURA = "01111" THEN
		SHLL <= '1';
	END IF;
	IF LECTURA = "10000" THEN
		SUB <= '1';
	END IF;
	IF LECTURA = "10001" THEN
		DEC <= '1';
	END IF;
	IF LECTURA = "10001" THEN
		JMP <= '1';
	END IF;
	IF MODO = '0' THEN
	   MODE <= '0';
	END IF;
	IF MODO ='1' THEN
		MODE <= '1';
	END IF;
END PROCESS;
END ESTRUCTURAL;
