library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.all;
USE ieee.std_logic_unsigned.all;

ENTITY DECODER2 IS --74_LS_42 MODIFICADO 
PORT (
	ENABLE_DEC: IN STD_LOGIC;
	IND: IN STD_LOGIC_VECTOR(7 downto 0);
	OP1: OUT STD_LOGIC_VECTOR(2 downto 0);
	OP2: OUT STD_LOGIC_VECTOR (2 downto 0)
);
END DECODER2
ARCHITECTURE ESTRUCTURAL OF DECODER2 IS
BEGIN
PROCESS (ENABLE_DEC)
	IF IND(7 DOWNTO 5) = "000" THEN
		OP1 <= R1;
	END IF;
	IF IND(7 DOWNTO 5) = "001" THEN
		OP1 <= R2;
	END IF;
	IF IND(7 DOWNTO 5) = "010" THEN
		OP1 <= R3;
	END IF;
	IF IND(7 DOWNTO 5) = "011" THEN
		OP1 <= R4;
	END IF;
	IF IND(7 DOWNTO 5) = "100" THEN
		OP1 <= RAUX;
	END IF;
	IF IND(7 DOWNTO 5) = "101" THEN
		OP1 <= RAUX2
	END IF;
	IF IND(4 DOWNTO 2) = "000" THEN
		OP2 <= R1;
	END IF;
	IF IND(4 DOWNTO 2) = "001" THEN
		OP2 <= R2;
	END IF;
	IF IND(4 DOWNTO 2) = "010" THEN
		OP2 <= R3;
	END IF;
	IF IND(4 DOWNTO 2) = "011" THEN
		OP2 <= R4;
	END IF;
	IF IND(4 DOWNTO 2) = "100" THEN
		OP2 <= RAUX;
	END IF;
	IF IND(4 DOWNTO 2) = "101" THEN
		OP2 <= RAUX2;
	END IF;
END PROCESS;
END ESTRUCTURAL;